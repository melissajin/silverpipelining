
module hazard_detection
(
    /* inputs */
    input logic i_mem_resp, d_mem_resp, d_mem_read,
    input lc3b_opcode op_MEM, op_WB,

    /* outputs */
    

);



endmodule // hazard_detection
