import lc3b_types::*;

module hardware_prefetcher
(

);

hardware_prefetcher_controller controller
(

);

hardware_prefetcher_datapath datapath
(

);


endmodule : hardware_prefetcher
