import lc3b_types::*;

module hardware_prefetcher_datapath
(

);

endmodule : hardware_prefetcher_datapath
