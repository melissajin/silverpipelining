import lc3b_types::*;

module ir_id_reg
(
    input clk,
    input load,
    input clear,
    input lc3b_word in,
    output lc3b_opcode opcode,
    output lc3b_reg dest, src1, src2,
    output lc3b_ir_10_0 ir_10_0
);

lc3b_word data;

always_ff @(posedge clk)
begin
    if(clear == 1)
      begin
        data = 0;
      end

    if (load == 1)
    begin
        data = in;
    end
end

always_comb
begin
    opcode = lc3b_opcode'(data[15:12]);

    dest = data[11:9];
    src1 = data[8:6];
    src2 = data[2:0];
    ir_10_0 = data[10:0];
end

endmodule : ir_id_reg
