import lc3b_types::*;

module hardware_prefetcher_controller
(

);

endmodule : hardware_prefetcher_controller
